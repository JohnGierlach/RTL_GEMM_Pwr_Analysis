`timescale 1ps/1ps

module gemm_top(
    input iclk, irst
    output
);


endmodule